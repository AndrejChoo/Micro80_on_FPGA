//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Tue Feb  3 11:33:23 2026

module zrom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h00000000000FFFFF00000000000FFFFF00000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h000000FFFFFFFFFF000000FFFFFFFFFF000000FFFFF00000000000FFFFF00000;
defparam prom_inst_0.INIT_RAM_02 = 256'h000000008888EC800000000C22A2A2C0000000088AEC08800000000CEE6E6EC0;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000008CE888800000000008CEC8000000000008CEC8000000000008CEEEC0;
defparam prom_inst_0.INIT_RAM_04 = 256'h00000000000FFFFF00000000000FFFFF00000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h000000FFFFFFFFFF000000FFFFFFFFFF000000FFFFF00000000000FFFFF00000;
defparam prom_inst_0.INIT_RAM_06 = 256'h000000CCCCCCCCCC0000000008CC800000000000C86EC80000000000C86E6880;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000008C4C80000000000BBBBF00000000000000E00000000000000FF0000;
defparam prom_inst_0.INIT_RAM_08 = 256'h00000000CCECECC00000000000004660000000008088CC800000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000880000000006CC68C80000000006608C60000000000C8CCC8C0;
defparam prom_inst_0.INIT_RAM_0A = 256'h00000000088E8800000000000C8E8C000000000008CCC80000000000C80008C0;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000008C60000000008800000000000000000E00000000000088000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h00000000C66C66C000000000E00C66C000000000E888888000000000C666E6C0;
defparam prom_inst_0.INIT_RAM_0D = 256'h000000000008C6E000000000C66C008000000000C66C00E000000000ECECCCC0;
defparam prom_inst_0.INIT_RAM_0E = 256'h00000000880088000000000088008800000000008C6E66C000000000C66C66C0;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000808C66C000000000008C80000000000000E0E000000000006C808C60;
defparam prom_inst_0.INIT_RAM_10 = 256'h00000000C60006C000000000C66C66C00000000066E666C000000000C0E6E6C0;
defparam prom_inst_0.INIT_RAM_11 = 256'h00000000C66E06C000000000000800E000000000E00800E0000000008C666C80;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000066C8C66000000000C66666E000000000C88888C000000000666E6660;
defparam prom_inst_0.INIT_RAM_13 = 256'h00000000C66666C00000000066EE666000000000666EEE6000000000E0000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000000C66C06C00000000066C666C00000000ECE6666C00000000000C666C0;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000CE666660000000008C66666000000000C666666000000000888888E0;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000C00000C000000000E008C6E000000000888C66600000000066C8C660;
defparam prom_inst_0.INIT_RAM_17 = 256'h00000000E0000000000000000006C80000000000CCCCCCC00000000026C80000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000003F666666000000000C666C0E00000000066E666C000000000C66666C0;
defparam prom_inst_0.INIT_RAM_19 = 256'h00000000000000E00000000000C666C000000000E00800E000000001F66666E0;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000066C8C66000000000666EE66800000000666EE6600000000066C8C660;
defparam prom_inst_0.INIT_RAM_1B = 256'h00000000C66666C000000000666E666000000000666EEE6000000000666666E0;
defparam prom_inst_0.INIT_RAM_1C = 256'h00000000C60006C00000000000C666C00000000066E666E000000000666666E0;
defparam prom_inst_0.INIT_RAM_1D = 256'h00000000C66C66C00000000066C8C66000000000C66E666000000000888888E0;
defparam prom_inst_0.INIT_RAM_1E = 256'h00000000E666666000000000C66C66C0000000006EEE666000000000C666C000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00000000EEEEEEE00000000066E6666000000003F666666000000000C66E66C0;
defparam prom_inst_0.INIT_RAM_20 = 256'h000000888888000000000088888F0000000000888888888800000000000F0000;
defparam prom_inst_0.INIT_RAM_21 = 256'h000000888888888800000088888F8888000000000008888800000000000F8888;
defparam prom_inst_0.INIT_RAM_22 = 256'h000000008CCCAEE000000088888F888800000000000F888800000088888F0000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000006CEC600000000000EE6E6E0000000000000E6E0000000000C08CC80;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000008CEC800000000D7D7D7D7D7000000A5A5A5A5A50000002828282828;
defparam prom_inst_0.INIT_RAM_25 = 256'h00000000C6C66C0C00000000AAAAAAE0000000008CE8EC8000000004CCCCCCC4;
defparam prom_inst_0.INIT_RAM_26 = 256'h00000000E00000000000000E8CE8EC8000000000EEE000000000000060666660;
defparam prom_inst_0.INIT_RAM_27 = 256'h00000000C66C000000000000088CCEE000000000EECC88000000000008CEC800;
defparam prom_inst_0.INIT_RAM_28 = 256'h00000000C0E6C0C00000008888F8F00000000066666666660000000000F0F000;
defparam prom_inst_0.INIT_RAM_29 = 256'h00000066666E00000000008888888000000000666670F00000000066666F0000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000000000F0766600000000000F66660000000000F8F888000000666666E000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000008888F8F8880000000000E6666600000000000E66660000000000888888;
defparam prom_inst_0.INIT_RAM_2C = 256'h00000000E00800EC000000888888888800000066667076660000006666676666;
defparam prom_inst_0.INIT_RAM_2D = 256'h00000066666F00000000008888F0F00000000066666666660000006666666666;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000F0766600000000000F66660000000000F0F888000000666670F000;
defparam prom_inst_0.INIT_RAM_2F = 256'h00000000C2A2A2C0000000666670766600000066666766660000008888F0F888;
defparam prom_inst_0.INIT_RAM_30 = 256'h00000000C606C00000000000C666C000000000006CCC8000000000000000C800;
defparam prom_inst_0.INIT_RAM_31 = 256'h00000008CCCC600000000000000806C000000000C0E6C000000000006CCCCCC0;
defparam prom_inst_0.INIT_RAM_32 = 256'h000000006C8C60000000000C6666606000000000C8888080000000006666C000;
defparam prom_inst_0.INIT_RAM_33 = 256'h00000000C666C000000000006666C00000000000666EC00000000000C8888880;
defparam prom_inst_0.INIT_RAM_34 = 256'h00000000C6C0E000000000000006C0000000000ECCCC6000000000000C66C000;
defparam prom_inst_0.INIT_RAM_35 = 256'h00000000CE666000000000008C666000000000006CCCC00000000000C600C000;
defparam prom_inst_0.INIT_RAM_36 = 256'h00000000E88088E000000000E08CE0000000000C6E666000000000006C8C6000;
defparam prom_inst_0.INIT_RAM_37 = 256'h00000000C6C000000000000000000C6000000000088E88000000000088808880;
defparam prom_inst_0.INIT_RAM_38 = 256'h00000006ECCCC00000000000C66C0C00000000006CCC800000000000C666C000;
defparam prom_inst_0.INIT_RAM_39 = 256'h000000000000E000000000000C66C00000000000C0E6C00000000006ECCCC000;
defparam prom_inst_0.INIT_RAM_3A = 256'h000000006C8C60000000000066EE68000000000066EE6000000000006C8C6000;
defparam prom_inst_0.INIT_RAM_3B = 256'h00000000C666C0000000000066E660000000000066EE6000000000006666E000;
defparam prom_inst_0.INIT_RAM_3C = 256'h00000000C606C0000000000000C6C0000000000066E6E000000000006666E000;
defparam prom_inst_0.INIT_RAM_3D = 256'h00000000C6C6C000000000006C8C600000000000C6E66000000000008888E000;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000E666600000000000C6C6C000000000006E66600000000000C6C00000;
defparam prom_inst_0.INIT_RAM_3F = 256'h00000000E66C80000000000066E6600000000003F666600000000000C6E6C000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h00000000000FFFFF000000000000000000000000000FFFFF0000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h00000000000FFFFF000000000000000000000000000FFFFF0000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h00000000111173100000000789B8A870000000022BF7133000000007FECFDF70;
defparam prom_inst_1.INIT_RAM_03 = 256'h000000001371111000000000010F010000000000137F731000000000137FFF60;
defparam prom_inst_1.INIT_RAM_04 = 256'h000000FFFFFFFFFF000000FFFFF00000000000FFFFFFFFFF000000FFFFF00000;
defparam prom_inst_1.INIT_RAM_05 = 256'h000000FFFFFFFFFF000000FFFFF00000000000FFFFFFFFFF000000FFFFF00000;
defparam prom_inst_1.INIT_RAM_06 = 256'h000000111111111100000000013310000000000073DF73100000000073DFD330;
defparam prom_inst_1.INIT_RAM_07 = 256'h000000000364630000000000117DDC7000000000036F63000000000000FF0000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000066F6F660000000000000266000000000101133100000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000003110000000007CD7363000000000C631CC0000000000C7CCC7C0;
defparam prom_inst_1.INIT_RAM_0A = 256'h000000000117110000000000063F360000000000310001300000000001333100;
defparam prom_inst_1.INIT_RAM_0B = 256'h000000008C631000000000001100000000000000000700000000000311000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h000000007C010C7000000000FC710C700000000071111310000000007CEDCC70;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000033310CF0000000007CCFC630000000007C0FCCF00000000010FC6310;
defparam prom_inst_1.INIT_RAM_0E = 256'h00000003110011000000000011001100000000007007CC70000000007CC7CC70;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000000010100C70000000006310136000000000007070000000000000131000;
defparam prom_inst_1.INIT_RAM_10 = 256'h000000007CCCCC7000000000FCCFCCF000000000CCFCCC70000000007CDDDC70;
defparam prom_inst_1.INIT_RAM_11 = 256'h000000007CCDCC7000000000CCCFCCF000000000FCCFCCF000000000FCCCCCF0;
defparam prom_inst_1.INIT_RAM_12 = 256'h00000000CCCFCCC0000000007CC00010000000003111113000000000CCCFCCC0;
defparam prom_inst_1.INIT_RAM_13 = 256'h000000007CCCCC7000000000CCCDFEC000000000CCDFFEC000000000FCCCCCC0;
defparam prom_inst_1.INIT_RAM_14 = 256'h000000007C07CC7000000000CCFCCCF0000000007CCCCC7000000000CCFCCCF0;
defparam prom_inst_1.INIT_RAM_15 = 256'h000000006FDDCCC00000000036CCCCC0000000007CCCCCC00000000011111170;
defparam prom_inst_1.INIT_RAM_16 = 256'h000000003333333000000000F63100F0000000001113666000000000CC636CC0;
defparam prom_inst_1.INIT_RAM_17 = 256'h00000000F000000000000000000C6310000000003000003000000000000136C0;
defparam prom_inst_1.INIT_RAM_18 = 256'h00000000FCCCCCC000000000FCCCFCF000000000CCFCCC7000000000DDDFDDD0;
defparam prom_inst_1.INIT_RAM_19 = 256'h00000000CCCCCCF000000000117DDD7000000000FCCFCCF00000000CF6666310;
defparam prom_inst_1.INIT_RAM_1A = 256'h00000000CCCFCCC000000000CEFDCCD300000000CEFDCCC000000000CC636CC0;
defparam prom_inst_1.INIT_RAM_1B = 256'h000000007CCCCC7000000000CCCFCCC000000000CCDFFEC000000000C6666310;
defparam prom_inst_1.INIT_RAM_1C = 256'h000000007CCCCC7000000000CCFCCCF000000000C67CCC7000000000CCCCCCF0;
defparam prom_inst_1.INIT_RAM_1D = 256'h00000000FCCFCCF000000000DD737DD0000000007C07CCC00000000011111170;
defparam prom_inst_1.INIT_RAM_1E = 256'h00000000FDDDDDD0000000007C010C7000000000FDDDFCC000000000FCCCFCC0;
defparam prom_inst_1.INIT_RAM_1F = 256'h00000000FFFFFFF000000000007CCCC000000000FDDDDDD0000000007C030C70;
defparam prom_inst_1.INIT_RAM_20 = 256'h00000011111F00000000001111110000000000111111111100000000000F0000;
defparam prom_inst_1.INIT_RAM_21 = 256'h00000011111F1111000000111111111100000000000F11110000000000011111;
defparam prom_inst_1.INIT_RAM_22 = 256'h000000007CCC701000000011111F111100000000000F111100000011111F0000;
defparam prom_inst_1.INIT_RAM_23 = 256'h000000001D7E7D1000000000EE66767000000000EF733330000000003F37CC70;
defparam prom_inst_1.INIT_RAM_24 = 256'h0000000233333332000000D7D7D7D7D7000000A5A5A5A5A50000002828282828;
defparam prom_inst_1.INIT_RAM_25 = 256'h000000003036636300000000117DDD7000000000137173100000000001373100;
defparam prom_inst_1.INIT_RAM_26 = 256'h00000000FCC00000000000071371731000000000777000000000000060666660;
defparam prom_inst_1.INIT_RAM_27 = 256'h00000000333333F00000000013377FF000000000FF77331000000000026F6200;
defparam prom_inst_1.INIT_RAM_28 = 256'h000000007CFC7060000000111111100000000033333333330000000000F0F000;
defparam prom_inst_1.INIT_RAM_29 = 256'h00000033333F00000000001111F1F00000000033333330000000003333330000;
defparam prom_inst_1.INIT_RAM_2A = 256'h0000000000333333000000000003333300000000001111110000003333F0F000;
defparam prom_inst_1.INIT_RAM_2B = 256'h00000011111111110000000000F0F33300000000000F33330000000000F1F111;
defparam prom_inst_1.INIT_RAM_2C = 256'h00000000FCCFCCF60000001111F1F11100000033333333330000003333333333;
defparam prom_inst_1.INIT_RAM_2D = 256'h00000033333F00000000001111F0F0000000003333F0F33300000033333F3333;
defparam prom_inst_1.INIT_RAM_2E = 256'h0000000000F0F33300000000000F33330000000000F0F1110000003333F0F000;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000078BAB8700000003333F0F33300000033333F33330000001111F0F111;
defparam prom_inst_1.INIT_RAM_30 = 256'h000000007CCC700000000000D66676E0000000007C7070000000000000000130;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000F07CC700000000000F66F6630000000007CFC7000000000007CCC7010;
defparam prom_inst_1.INIT_RAM_32 = 256'h00000000E67666E00000000366000000000000003111301000000000E66766E0;
defparam prom_inst_1.INIT_RAM_33 = 256'h000000007CCC7000000000006666D00000000000DDDFE0000000000031111130;
defparam prom_inst_1.INIT_RAM_34 = 256'h00000000F07C700000000000F667D0000000000107CC70000000000F6766D000;
defparam prom_inst_1.INIT_RAM_35 = 256'h000000006FDDC0000000000036CCC000000000007CCCC000000000001333F330;
defparam prom_inst_1.INIT_RAM_36 = 256'h000000000117110000000000731070000000000707CCC00000000000C636C000;
defparam prom_inst_1.INIT_RAM_37 = 256'h000000003333F0000000000000000D7000000000711011700000000011101110;
defparam prom_inst_1.INIT_RAM_38 = 256'h00000000FCCCC000000000007CC7C700000000007C70700000000000DDFDD000;
defparam prom_inst_1.INIT_RAM_39 = 256'h00000000CCCCF0000000000017DD7000000000007CFC70000000000CF6663000;
defparam prom_inst_1.INIT_RAM_3A = 256'h00000000E676E00000000000EFDCC30000000000EFDCC00000000000C636C000;
defparam prom_inst_1.INIT_RAM_3B = 256'h000000007CCC700000000000CCFCC00000000000CDFEC00000000000E6663000;
defparam prom_inst_1.INIT_RAM_3C = 256'h000000007CCC7000000000006676700000000000C67C700000000000CCCCF000;
defparam prom_inst_1.INIT_RAM_3D = 256'h00000000FCFCF00000000000D737D00000000000707CC0000000000011117000;
defparam prom_inst_1.INIT_RAM_3E = 256'h00000000FDDDD000000000007C1C700000000000FDFCC00000000000FCFCC000;
defparam prom_inst_1.INIT_RAM_3F = 256'h00000000FCC6310000000000007CC00000000000FDDDD000000000007C1C7000;

endmodule //zrom
